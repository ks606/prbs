/********************************************************************************/
// Engineer:        
// Design Name: PRBS_TX
// Module Name: PRBS_TX     
// Target Device:    
// Description: PRBS transceiver
//      
// Dependencies:
//    None
// Revision:
//    None
// Additional Comments: 
//
/********************************************************************************/

`ifndef _PRBS_TX
`define _PRBS_TX

module PRBS_TX #(parameter 
							PRBS_TYPE = 7

)(
	input 					clk,
	input 					rst,
	
	// Input interface
	input 					prbs_en,
	
	// Output interface
	output 					dout_vld,
	output 					dout
	
);

/********************************************************************************/
// Parameters section
/********************************************************************************/ 
/********************************************************************************/
// Signals declaration section
/********************************************************************************/


/********************************************************************************/
// Main section
/********************************************************************************/	
	wire [31:0]				gen_shift_reg;
	
	PRBS_GEN #(
        .PRBS_TYPE(PRBS_TYPE)
    )_PRBS_GEN(
        .clk				(clk), 
		.rst				(rst),
		// Input
		.prbs_en			(prbs_en), 
        
        // Output
		.gen_shift_reg		(gen_shift_reg),
        .dout				(dout),
		.dout_vld			(dout_vld)
	
	);
	
	/****************************************************************************/
    // Delay
    /****************************************************************************/  

	
	/****************************************************************************/
    // Input bit counter
    /****************************************************************************/ 

	
	/****************************************************************************/
    // Shift register
    /****************************************************************************/ 

	/****************************************************************************/
    // Frame register
    /****************************************************************************/ 

	/****************************************************************************/
    // 
    /****************************************************************************/	
		
		
	
	/****************************************************************************/
    // Error/data counters
    /****************************************************************************/ 	


/********************************************************************************/
// Output
/********************************************************************************/

	
endmodule

`endif // _PRBS_TX